VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO LOGIC0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LOGIC0 0 0 ;
  SIZE 175 BY 1402 ;
  SYMMETRY X Y ;
  SITE std_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal2 ;
        RECT 0 1320 630 1470 ;
        RECT 175 275 225 1470 ;
        RECT 100 275 150 1470 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal2 ;
        RECT 0 0 630 150 ;
        RECT 555 0 605 1195 ;
    END
  END VSS
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 36.25 1065 141.25 1170 ;
    END
  END OUT
  PIN VBG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0 150 175 200 ;
        RECT 0 1270 175 1320 ;
    END
  END VBG
  OBS
    LAYER metal2 ;
      RECT 36.25 1065 141.25 1170 ;
      RECT 38.4 0 138.4 1170 ;
      RECT 37 1401 40.5 1402 ;
      RECT 41 1396 42 1401 ;
      RECT 40 1400.75 42 1401 ;
      RECT 40.5 1400.25 41 1401.75 ;
      RECT 37 1395 38 1402 ;
      RECT 40.5 1395.25 41 1396.75 ;
      RECT 40 1396 42 1396.25 ;
      RECT 37 1395 40.5 1396 ;
      RECT 31 1401 34.5 1402 ;
      RECT 35 1396 36 1401 ;
      RECT 34 1400.75 36 1401 ;
      RECT 34.5 1400.25 35 1401.75 ;
      RECT 31 1395 32 1402 ;
      RECT 34.5 1395.25 35 1396.75 ;
      RECT 34 1396 36 1396.25 ;
      RECT 31 1395 34.5 1396 ;
      RECT 29 1396.5 30 1402 ;
      RECT 25 1396.5 26 1402 ;
      RECT 28 1395.5 29 1397 ;
      RECT 26 1395.5 27 1397 ;
      RECT 27 1395 28 1396.25 ;
  END
END LOGIC0

END LIBRARY
